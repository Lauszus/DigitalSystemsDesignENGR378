library verilog;
use verilog.vl_types.all;
entity t_two_bit_counter is
end t_two_bit_counter;
