library verilog;
use verilog.vl_types.all;
entity t_JK is
end t_JK;
